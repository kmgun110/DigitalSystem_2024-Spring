library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Full_Adder is
    port(x, y, cin : in std_logic; -- entity�� input�� x, y, cin
    sum : out std_logic;
    cout : out std_logic);  -- entity�� output�� sum, cout
end Full_Adder;

architecture Behavioral of Full_Adder is

begin -- Full Adder���� sum�� cout�� ���� 
    sum <= cin xor (x xor y);
    cout <= (x and y) or (x and cin) or (y and cin);

end Behavioral;
