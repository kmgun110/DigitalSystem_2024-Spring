library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Adder_4bit is
    port (x, y: in std_logic_vector(3 downto 0);   -- entity�� input�� x, y, cin
    cin : in std_logic;                             -- �� ��, x, y�� 4-bit vector
    sum : out std_logic_vector(3 downto 0);   -- entity�� output�� sum, cout
    cout : out std_logic);                     -- �� ��, sum�� 4-bit vector
end Adder_4bit;

architecture Behavioral of Adder_4bit is
component Full_Adder   -- Full_Adder�� component�� �ҷ���
    port (x, y, cin : in std_logic;
    sum, cout : out std_logic);
end component;

signal c : std_logic_vector(3 downto 1);   -- �� Full Adder�� cout�� bit vector�� ����

begin
    FA0: Full_Adder port map(x(0), y(0), cin, sum(0), c(1));   -- ù��° Full Adder
    FA1: Full_Adder port map(x(1), y(1), c(1), sum(1), c(2));   -- �ι�° Full Adder
    FA2: Full_Adder port map(x(2), y(2), c(2), sum(2), c(3));   -- ����° Full Adder
    FA3: Full_Adder port map(x(3), y(3), c(3), sum(3), cout);   -- �׹�° Full Adder
end Behavioral;
