library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Full_Adder_tb is
end Full_Adder_tb;

architecture Behavioral of Full_Adder_tb is
    component Full_Adder port(  -- �ռ� ������ Full_Adder�� component �ҷ���
        x, y, cin : in std_logic;
        sum : out std_logic;
        cout : out std_logic); 
    end component;   
    
    signal X : std_logic :='0';   -- X, Y, Cin�� �ʱⰪ ����
    signal Y : std_logic :='1';
    signal Cin : std_logic :='1';
    signal Sum, Cout : std_logic; 
    
begin
    uut : Full_Adder port map (
        x => X,   -- �ҷ��� Full_Adder�� component�� ������ signal�� �Ҵ�
        y => Y,
        cin => Cin,
        sum => Sum,
        cout => Cout);
stim_proc : process
    begin
    X <= '1'; 
    Y <= '1';  
    wait for 10ns;  
    Cin <= '0';  -- 10ns ���� Cin = 0
    wait for 10ns;
    X <= '0';  -- 10ns ���� X = 0, Y = 0, Cin = 1
    Y <= '0';
    Cin <= '1';
    wait for 10ns;
    Cin <= '0';   -- 10ns ���� Cin = 0
    wait for 10ns;
    X <= '1';   -- 10ns ���� X = 1, Y =1 0
    Y <= '0';
    wait for 10ns;   -- 10ns ���� process���� ó������ ���ư�
  end process;
  
end Behavioral;
